.SUBCKT PSRMINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=450n L=60n M=1
.ENDS

.SUBCKT PSRMBUF A Z VDD VSS
MPM0 n1 A VDD VDD P_12_LLRVT W=210n L=60n M=1
MNM0 n1 A VSS VSS N_12_LLRVT W=150n L=60n M=1
MPM1 Z n1 VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM1 Z n1 VSS VSS N_12_LLRVT W=450n L=60n M=1
.ENDS

.SUBCKT PSRMND A B Z VDD VSS
*.PININFO A:I B:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=270n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=270n L=60n M=1
MNM0 Z B n1 VSS N_12_LLRVT W=180n L=60n M=1
MNM1 n1 A VSS VSS N_12_LLRVT W=180n L=60n M=1
.ENDS

.SUBCKT PSRMNR A B Z VDD VSS
*.PININFO A:I B:I Z:O
MPM0 n1 A VDD VDD P_12_LLRVT W=270n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=270n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=180n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=180n L=60n M=1
.ENDS

.SUBCKT PSADOH_ND2 A B Z VDD VSS
*.PININFO A:I B:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z B n1 VSS N_12_LLRVT W=480n L=60n M=1
MNM1 n1 A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_ND3 A B C Z VDD VSS
*.PININFO A:I B:I C:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM2 Z C VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z C n1 VSS N_12_LLRVT W=480n L=60n M=1
MNM1 n1 B n2 VSS N_12_LLRVT W=480n L=60n M=1
MNM2 n2 A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_NR2 A B Z VDD VSS
*.PININFO A:I B:I Z:O
MPM0 n1 A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_NR3 A B C Z VDD VSS
*.PININFO A:I B:I C:I Z:O VDD:B VSS:B
MPM0 Z  C n1  VDD P_12_LLRVT W=660n L=60n M=1
MPM1 n1 B n2  VDD P_12_LLRVT W=660n L=60n M=1
MPM2 n2 A VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z  A VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM1 Z  B VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM2 Z  C VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSREG_LA1 D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSREG_LA2 D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=300n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=450n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSREG D CKP CKN QP QN VDD VSS
XI0 D CKN CKP n1 i1 VDD VSS PSREG_LA1
XI1 n1 CKP CKN QP QN VDD VSS PSREG_LA2
.ENDS

.SUBCKT PSADCKG_LA D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSADCKG_NR2 A B Z VDD VSS
MPM0 n1 A VDD VDD P_12_LLRVT W=630n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSADCKG E CKP CKN GCKP GCKN VDD VSS
X1 E CKN CKP i1 n1 VDD VSS PSADCKG_LA
X2 n1 CKN n2 VDD VSS PSADCKG_NR2
MPM0 GCKN n2 VDD VDD P_12_LLRVT W=600n L=60n M=1
MNM0 GCKN n2 VSS VSS N_12_LLRVT W=300n L=60n M=1
MPM1 GCKP GCKN VDD VDD P_12_LLRVT W=600n L=60n M=1
MNM1 GCKP GCKN VSS VSS N_12_LLRVT W=300n L=60n M=1
.ENDS

.SUBCKT PSADINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSBA1 D GP GN S Q VDD VSS
*.PININFO D:I GP:I GN:I S:I Q:O VDD:B VSS:B
MNM0 net41 D VSS VSS N_12_LLRVT W=200e-9 L=60n M=1
MNM1 nFB GP net41 VSS N_12_LLRVT W=200e-9 L=60n M=1
MNM2 net40 nZ VSS VSS N_12_LLRVT W=150e-9 L=60n M=1
MNM3 nFB GN net40 VSS N_12_LLRVT W=150e-9 L=60n M=1
MNM4 nZ nFB VSS VSS N_12_LLRVT W=180e-9 L=60n M=1
MNM5 net42 S VSS VSS N_12_LLRVT W=180e-9 L=60n M=1
MNM6 Q nZ net42 VSS N_12_LLRVT W=180e-9 L=60n M=1
MPM0 nFB GN net38 VDD P_12_LLRVT W=300e-9 L=60n M=1
MPM1 net38 D VDD VDD P_12_LLRVT W=300e-9 L=60n M=1
MPM2 nFB GP net39 VDD P_12_LLRVT W=150e-9 L=60n M=1
MPM3 net39 nZ VDD VDD P_12_LLRVT W=150e-9 L=60n M=1
MPM4 nZ nFB VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
MPM5 Q nZ VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
MPM6 Q S VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
.ENDS

.SUBCKT PSRWCKG_CKINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=260n L=60n M=1
.ENDS

.SUBCKT PSRWCKG RE WE CK RCKP RCKN WCKP WCKN VDD VSS
X0 RE nCKP nCKN RCKP RCKN VDD VSS PSADCKG
X1 WE nCKP nCKN WCKP WCKN VDD VSS PSADCKG
X2 CK nCKN VDD VSS PSRWCKG_CKINV
X3 nCKN nCKP VDD VSS PSRWCKG_CKINV
.ENDS


.SUBCKT PSADOH4R A0 A1 Z VDD VSS
*.PININFO A0:I A1:I Z:O VDD:B VSS:B
X0 A0 A1 Z VDD VSS PSADOH_NR2
.ENDS

.SUBCKT PSADOH4 A0 A1 Z0 Z1 Z2 Z3 VDD VSS
XI0 A0 N0 VDD VSS PSADINV
XI1 A1 N1 VDD VSS PSADINV
X0 A0 A1 Z0 VDD VSS PSADOH4R
X1 N0 A1 Z1 VDD VSS PSADOH4R
X2 A0 N1 Z2 VDD VSS PSADOH4R
X3 N0 N1 Z3 VDD VSS PSADOH4R
.ENDS

.SUBCKT PSAD4 CKP CKN RA0 RA1 WA0 WA1 S0 GP0 GN0 S1 GP1 GN1 S2 GP2 GN2 S3 GP3 GN3 VDD VSS
XCKG0 nWE0 CKP CKN GP0 GN0 VDD VSS PSADCKG 
XCKG1 nWE1 CKP CKN GP1 GN1 VDD VSS PSADCKG 
XCKG2 nWE2 CKP CKN GP2 GN2 VDD VSS PSADCKG 
XCKG3 nWE3 CKP CKN GP3 GN3 VDD VSS PSADCKG 
XRAD RA0 RA1 S0 S1 S2 S3 VDD VSS PSADOH4
XWAD WA0 WA1 nWE0 nWE1 nWE2 nWE3 VDD VSS PSADOH4
.ENDS

.SUBCKT PSBA4 D S0 GP0 GN0 S1 GP1 GN1 S2 GP2 GN2 S3 GP3 GN3 Q VDD VSS
X0 D GP0 GN0 S0 nL0Q0 VDD VSS PSBA1
X1 D GP1 GN1 S1 nL0Q1 VDD VSS PSBA1
X2 D GP2 GN2 S2 nL0Q2 VDD VSS PSBA1
X3 D GP3 GN3 S3 nL0Q3 VDD VSS PSBA1
XINV nQ Q VDD VSS PSRMINV
XL1Q0 nL0Q0 nL0Q1 nL1Q0 VDD VSS PSRMND
XL1Q1 nL0Q2 nL0Q3 nL1Q1 VDD VSS PSRMND
XL2Q0 nL1Q0 nL1Q1 nQ VDD VSS PSRMNR
.ENDS

.SUBCKT PS4X8 CK RE RA0 RA1 RD0 RD1 RD2 RD3 RD4 RD5 RD6 RD7 WE WA0 WA1 WD0 WD1 WD2 WD3 WD4 WD5 WD6 WD7 VDD VSS
XRWCKG RE WE CK nRCKP nRCKN nWCKP nWCKN VDD VSS PSRWCKG
XAD nWCKP nWCKN nRA0 nRA1 WA0 WA1 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 VDD VSS PSAD4
XWDREG0 WD0 nWCKP nWCKN nWD0 iw0 VDD VSS PSREG
XWDREG1 WD1 nWCKP nWCKN nWD1 iw1 VDD VSS PSREG
XWDREG2 WD2 nWCKP nWCKN nWD2 iw2 VDD VSS PSREG
XWDREG3 WD3 nWCKP nWCKN nWD3 iw3 VDD VSS PSREG
XWDREG4 WD4 nWCKP nWCKN nWD4 iw4 VDD VSS PSREG
XWDREG5 WD5 nWCKP nWCKN nWD5 iw5 VDD VSS PSREG
XWDREG6 WD6 nWCKP nWCKN nWD6 iw6 VDD VSS PSREG
XWDREG7 WD7 nWCKP nWCKN nWD7 iw7 VDD VSS PSREG
XRAREG0 RA0 nRCKP nRCKN nRA0 ir0 VDD VSS PSREG
XRAREG1 RA1 nRCKP nRCKN nRA1 ir1 VDD VSS PSREG
XBA0 nWD0 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD0 VDD VSS PSBA4
XBA1 nWD1 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD1 VDD VSS PSBA4
XBA2 nWD2 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD2 VDD VSS PSBA4
XBA3 nWD3 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD3 VDD VSS PSBA4
XBA4 nWD4 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD4 VDD VSS PSBA4
XBA5 nWD5 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD5 VDD VSS PSBA4
XBA6 nWD6 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD6 VDD VSS PSBA4
XBA7 nWD7 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD7 VDD VSS PSBA4
.ENDS
