.SUBCKT PSRMINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=450n L=60n M=1
.ENDS

.SUBCKT PSRMBUF A Z VDD VSS
MPM0 n1 A VDD VDD P_12_LLRVT W=210n L=60n M=1
MNM0 n1 A VSS VSS N_12_LLRVT W=150n L=60n M=1
MPM1 Z n1 VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM1 Z n1 VSS VSS N_12_LLRVT W=450n L=60n M=1
.ENDS

.SUBCKT PSRMND A B Z VDD VSS
*.PININFO A:I B:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=270n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=270n L=60n M=1
MNM0 Z B n1 VSS N_12_LLRVT W=180n L=60n M=1
MNM1 n1 A VSS VSS N_12_LLRVT W=180n L=60n M=1
.ENDS

.SUBCKT PSRMNR A B Z VDD VSS
*.PININFO A:I B:I Z:O
MPM0 n1 A VDD VDD P_12_LLRVT W=270n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=270n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=180n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=180n L=60n M=1
.ENDS

.SUBCKT PSADOH_ND2 A B Z VDD VSS
*.PININFO A:I B:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z B n1 VSS N_12_LLRVT W=480n L=60n M=1
MNM1 n1 A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_ND3 A B C Z VDD VSS
*.PININFO A:I B:I C:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM2 Z C VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z C n1 VSS N_12_LLRVT W=480n L=60n M=1
MNM1 n1 B n2 VSS N_12_LLRVT W=480n L=60n M=1
MNM2 n2 A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_NR2 A B Z VDD VSS
*.PININFO A:I B:I Z:O
MPM0 n1 A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_NR3 A B C Z VDD VSS
*.PININFO A:I B:I C:I Z:O VDD:B VSS:B
MPM0 Z  C n1  VDD P_12_LLRVT W=660n L=60n M=1
MPM1 n1 B n2  VDD P_12_LLRVT W=660n L=60n M=1
MPM2 n2 A VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z  A VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM1 Z  B VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM2 Z  C VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSREG_LA1 D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSREG_LA2 D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=300n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=450n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSREG D CKP CKN QP QN VDD VSS
XI0 D CKN CKP n1 i1 VDD VSS PSREG_LA1
XI1 n1 CKP CKN QP QN VDD VSS PSREG_LA2
.ENDS

.SUBCKT PSADCKG_LA D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSADCKG_NR2 A B Z VDD VSS
MPM0 n1 A VDD VDD P_12_LLRVT W=630n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSADCKG E CKP CKN GCKP GCKN VDD VSS
X1 E CKN CKP i1 n1 VDD VSS PSADCKG_LA
X2 n1 CKN n2 VDD VSS PSADCKG_NR2
MPM0 GCKN n2 VDD VDD P_12_LLRVT W=600n L=60n M=1
MNM0 GCKN n2 VSS VSS N_12_LLRVT W=300n L=60n M=1
MPM1 GCKP GCKN VDD VDD P_12_LLRVT W=600n L=60n M=1
MNM1 GCKP GCKN VSS VSS N_12_LLRVT W=300n L=60n M=1
.ENDS

.SUBCKT PSADINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSBA1 D GP GN S Q VDD VSS
*.PININFO D:I GP:I GN:I S:I Q:O VDD:B VSS:B
MNM0 net41 D VSS VSS N_12_LLRVT W=200e-9 L=60n M=1
MNM1 nFB GP net41 VSS N_12_LLRVT W=200e-9 L=60n M=1
MNM2 net40 nZ VSS VSS N_12_LLRVT W=150e-9 L=60n M=1
MNM3 nFB GN net40 VSS N_12_LLRVT W=150e-9 L=60n M=1
MNM4 nZ nFB VSS VSS N_12_LLRVT W=180e-9 L=60n M=1
MNM5 net42 S VSS VSS N_12_LLRVT W=180e-9 L=60n M=1
MNM6 Q nZ net42 VSS N_12_LLRVT W=180e-9 L=60n M=1
MPM0 nFB GN net38 VDD P_12_LLRVT W=300e-9 L=60n M=1
MPM1 net38 D VDD VDD P_12_LLRVT W=300e-9 L=60n M=1
MPM2 nFB GP net39 VDD P_12_LLRVT W=150e-9 L=60n M=1
MPM3 net39 nZ VDD VDD P_12_LLRVT W=150e-9 L=60n M=1
MPM4 nZ nFB VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
MPM5 Q nZ VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
MPM6 Q S VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
.ENDS

.SUBCKT PSRWCKG_CKINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=260n L=60n M=1
.ENDS

.SUBCKT PSRWCKG RE WE CK RCKP RCKN WCKP WCKN VDD VSS
X0 RE nCKP nCKN RCKP RCKN VDD VSS PSADCKG
X1 WE nCKP nCKN WCKP WCKN VDD VSS PSADCKG
X2 CK nCKN VDD VSS PSRWCKG_CKINV
X3 nCKN nCKP VDD VSS PSRWCKG_CKINV
.ENDS


.SUBCKT PSADOH32R A0 A1 A2 A3 A4 Z VDD VSS
*.PININFO A0:I A1:I A2:I A3:I A4:I Z:O VDD:B VSS:B
X0 A0 A1 n1 VDD VSS PSADOH_ND2
X1 A2 A3 A4 n2 VDD VSS PSADOH_ND3
X2 n1 n2 Z VDD VSS PSADOH_NR2
.ENDS

.SUBCKT PSADOH32 A0 A1 A2 A3 A4 Z0 Z1 Z2 Z3 Z4 Z5 Z6 Z7 Z8 Z9 Z10 Z11 Z12 Z13 Z14 Z15 Z16 Z17 Z18 Z19 Z20 Z21 Z22 Z23 Z24 Z25 Z26 Z27 Z28 Z29 Z30 Z31 VDD VSS
XI0 A0 N0 VDD VSS PSADINV
XI1 A1 N1 VDD VSS PSADINV
XI2 A2 N2 VDD VSS PSADINV
XI3 A3 N3 VDD VSS PSADINV
XI4 A4 N4 VDD VSS PSADINV
X0 N0 N1 N2 N3 N4 Z0 VDD VSS PSADOH32R
X1 A0 N1 N2 N3 N4 Z1 VDD VSS PSADOH32R
X2 N0 A1 N2 N3 N4 Z2 VDD VSS PSADOH32R
X3 A0 A1 N2 N3 N4 Z3 VDD VSS PSADOH32R
X4 N0 N1 A2 N3 N4 Z4 VDD VSS PSADOH32R
X5 A0 N1 A2 N3 N4 Z5 VDD VSS PSADOH32R
X6 N0 A1 A2 N3 N4 Z6 VDD VSS PSADOH32R
X7 A0 A1 A2 N3 N4 Z7 VDD VSS PSADOH32R
X8 N0 N1 N2 A3 N4 Z8 VDD VSS PSADOH32R
X9 A0 N1 N2 A3 N4 Z9 VDD VSS PSADOH32R
X10 N0 A1 N2 A3 N4 Z10 VDD VSS PSADOH32R
X11 A0 A1 N2 A3 N4 Z11 VDD VSS PSADOH32R
X12 N0 N1 A2 A3 N4 Z12 VDD VSS PSADOH32R
X13 A0 N1 A2 A3 N4 Z13 VDD VSS PSADOH32R
X14 N0 A1 A2 A3 N4 Z14 VDD VSS PSADOH32R
X15 A0 A1 A2 A3 N4 Z15 VDD VSS PSADOH32R
X16 N0 N1 N2 N3 A4 Z16 VDD VSS PSADOH32R
X17 A0 N1 N2 N3 A4 Z17 VDD VSS PSADOH32R
X18 N0 A1 N2 N3 A4 Z18 VDD VSS PSADOH32R
X19 A0 A1 N2 N3 A4 Z19 VDD VSS PSADOH32R
X20 N0 N1 A2 N3 A4 Z20 VDD VSS PSADOH32R
X21 A0 N1 A2 N3 A4 Z21 VDD VSS PSADOH32R
X22 N0 A1 A2 N3 A4 Z22 VDD VSS PSADOH32R
X23 A0 A1 A2 N3 A4 Z23 VDD VSS PSADOH32R
X24 N0 N1 N2 A3 A4 Z24 VDD VSS PSADOH32R
X25 A0 N1 N2 A3 A4 Z25 VDD VSS PSADOH32R
X26 N0 A1 N2 A3 A4 Z26 VDD VSS PSADOH32R
X27 A0 A1 N2 A3 A4 Z27 VDD VSS PSADOH32R
X28 N0 N1 A2 A3 A4 Z28 VDD VSS PSADOH32R
X29 A0 N1 A2 A3 A4 Z29 VDD VSS PSADOH32R
X30 N0 A1 A2 A3 A4 Z30 VDD VSS PSADOH32R
X31 A0 A1 A2 A3 A4 Z31 VDD VSS PSADOH32R
.ENDS

.SUBCKT PSAD32 CKP CKN RA0 RA1 RA2 RA3 RA4 WA0 WA1 WA2 WA3 WA4 S0 GP0 GN0 S1 GP1 GN1 S2 GP2 GN2 S3 GP3 GN3 S4 GP4 GN4 S5 GP5 GN5 S6 GP6 GN6 S7 GP7 GN7 S8 GP8 GN8 S9 GP9 GN9 S10 GP10 GN10 S11 GP11 GN11 S12 GP12 GN12 S13 GP13 GN13 S14 GP14 GN14 S15 GP15 GN15 S16 GP16 GN16 S17 GP17 GN17 S18 GP18 GN18 S19 GP19 GN19 S20 GP20 GN20 S21 GP21 GN21 S22 GP22 GN22 S23 GP23 GN23 S24 GP24 GN24 S25 GP25 GN25 S26 GP26 GN26 S27 GP27 GN27 S28 GP28 GN28 S29 GP29 GN29 S30 GP30 GN30 S31 GP31 GN31 VDD VSS
XCKG0 nWE0 CKP CKN GP0 GN0 VDD VSS PSADCKG 
XCKG1 nWE1 CKP CKN GP1 GN1 VDD VSS PSADCKG 
XCKG2 nWE2 CKP CKN GP2 GN2 VDD VSS PSADCKG 
XCKG3 nWE3 CKP CKN GP3 GN3 VDD VSS PSADCKG 
XCKG4 nWE4 CKP CKN GP4 GN4 VDD VSS PSADCKG 
XCKG5 nWE5 CKP CKN GP5 GN5 VDD VSS PSADCKG 
XCKG6 nWE6 CKP CKN GP6 GN6 VDD VSS PSADCKG 
XCKG7 nWE7 CKP CKN GP7 GN7 VDD VSS PSADCKG 
XCKG8 nWE8 CKP CKN GP8 GN8 VDD VSS PSADCKG 
XCKG9 nWE9 CKP CKN GP9 GN9 VDD VSS PSADCKG 
XCKG10 nWE10 CKP CKN GP10 GN10 VDD VSS PSADCKG 
XCKG11 nWE11 CKP CKN GP11 GN11 VDD VSS PSADCKG 
XCKG12 nWE12 CKP CKN GP12 GN12 VDD VSS PSADCKG 
XCKG13 nWE13 CKP CKN GP13 GN13 VDD VSS PSADCKG 
XCKG14 nWE14 CKP CKN GP14 GN14 VDD VSS PSADCKG 
XCKG15 nWE15 CKP CKN GP15 GN15 VDD VSS PSADCKG 
XCKG16 nWE16 CKP CKN GP16 GN16 VDD VSS PSADCKG 
XCKG17 nWE17 CKP CKN GP17 GN17 VDD VSS PSADCKG 
XCKG18 nWE18 CKP CKN GP18 GN18 VDD VSS PSADCKG 
XCKG19 nWE19 CKP CKN GP19 GN19 VDD VSS PSADCKG 
XCKG20 nWE20 CKP CKN GP20 GN20 VDD VSS PSADCKG 
XCKG21 nWE21 CKP CKN GP21 GN21 VDD VSS PSADCKG 
XCKG22 nWE22 CKP CKN GP22 GN22 VDD VSS PSADCKG 
XCKG23 nWE23 CKP CKN GP23 GN23 VDD VSS PSADCKG 
XCKG24 nWE24 CKP CKN GP24 GN24 VDD VSS PSADCKG 
XCKG25 nWE25 CKP CKN GP25 GN25 VDD VSS PSADCKG 
XCKG26 nWE26 CKP CKN GP26 GN26 VDD VSS PSADCKG 
XCKG27 nWE27 CKP CKN GP27 GN27 VDD VSS PSADCKG 
XCKG28 nWE28 CKP CKN GP28 GN28 VDD VSS PSADCKG 
XCKG29 nWE29 CKP CKN GP29 GN29 VDD VSS PSADCKG 
XCKG30 nWE30 CKP CKN GP30 GN30 VDD VSS PSADCKG 
XCKG31 nWE31 CKP CKN GP31 GN31 VDD VSS PSADCKG 
XRAD RA0 RA1 RA2 RA3 RA4 S0 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13 S14 S15 S16 S17 S18 S19 S20 S21 S22 S23 S24 S25 S26 S27 S28 S29 S30 S31 VDD VSS PSADOH32
XWAD WA0 WA1 WA2 WA3 WA4 nWE0 nWE1 nWE2 nWE3 nWE4 nWE5 nWE6 nWE7 nWE8 nWE9 nWE10 nWE11 nWE12 nWE13 nWE14 nWE15 nWE16 nWE17 nWE18 nWE19 nWE20 nWE21 nWE22 nWE23 nWE24 nWE25 nWE26 nWE27 nWE28 nWE29 nWE30 nWE31 VDD VSS PSADOH32
.ENDS

.SUBCKT PSBA32 D S0 GP0 GN0 S1 GP1 GN1 S2 GP2 GN2 S3 GP3 GN3 S4 GP4 GN4 S5 GP5 GN5 S6 GP6 GN6 S7 GP7 GN7 S8 GP8 GN8 S9 GP9 GN9 S10 GP10 GN10 S11 GP11 GN11 S12 GP12 GN12 S13 GP13 GN13 S14 GP14 GN14 S15 GP15 GN15 S16 GP16 GN16 S17 GP17 GN17 S18 GP18 GN18 S19 GP19 GN19 S20 GP20 GN20 S21 GP21 GN21 S22 GP22 GN22 S23 GP23 GN23 S24 GP24 GN24 S25 GP25 GN25 S26 GP26 GN26 S27 GP27 GN27 S28 GP28 GN28 S29 GP29 GN29 S30 GP30 GN30 S31 GP31 GN31 Q VDD VSS
X0 D GP0 GN0 S0 nL0Q0 VDD VSS PSBA1
X1 D GP1 GN1 S1 nL0Q1 VDD VSS PSBA1
X2 D GP2 GN2 S2 nL0Q2 VDD VSS PSBA1
X3 D GP3 GN3 S3 nL0Q3 VDD VSS PSBA1
X4 D GP4 GN4 S4 nL0Q4 VDD VSS PSBA1
X5 D GP5 GN5 S5 nL0Q5 VDD VSS PSBA1
X6 D GP6 GN6 S6 nL0Q6 VDD VSS PSBA1
X7 D GP7 GN7 S7 nL0Q7 VDD VSS PSBA1
X8 D GP8 GN8 S8 nL0Q8 VDD VSS PSBA1
X9 D GP9 GN9 S9 nL0Q9 VDD VSS PSBA1
X10 D GP10 GN10 S10 nL0Q10 VDD VSS PSBA1
X11 D GP11 GN11 S11 nL0Q11 VDD VSS PSBA1
X12 D GP12 GN12 S12 nL0Q12 VDD VSS PSBA1
X13 D GP13 GN13 S13 nL0Q13 VDD VSS PSBA1
X14 D GP14 GN14 S14 nL0Q14 VDD VSS PSBA1
X15 D GP15 GN15 S15 nL0Q15 VDD VSS PSBA1
X16 D GP16 GN16 S16 nL0Q16 VDD VSS PSBA1
X17 D GP17 GN17 S17 nL0Q17 VDD VSS PSBA1
X18 D GP18 GN18 S18 nL0Q18 VDD VSS PSBA1
X19 D GP19 GN19 S19 nL0Q19 VDD VSS PSBA1
X20 D GP20 GN20 S20 nL0Q20 VDD VSS PSBA1
X21 D GP21 GN21 S21 nL0Q21 VDD VSS PSBA1
X22 D GP22 GN22 S22 nL0Q22 VDD VSS PSBA1
X23 D GP23 GN23 S23 nL0Q23 VDD VSS PSBA1
X24 D GP24 GN24 S24 nL0Q24 VDD VSS PSBA1
X25 D GP25 GN25 S25 nL0Q25 VDD VSS PSBA1
X26 D GP26 GN26 S26 nL0Q26 VDD VSS PSBA1
X27 D GP27 GN27 S27 nL0Q27 VDD VSS PSBA1
X28 D GP28 GN28 S28 nL0Q28 VDD VSS PSBA1
X29 D GP29 GN29 S29 nL0Q29 VDD VSS PSBA1
X30 D GP30 GN30 S30 nL0Q30 VDD VSS PSBA1
X31 D GP31 GN31 S31 nL0Q31 VDD VSS PSBA1
XBUF nQ Q VDD VSS PSRMBUF
XL1Q0 nL0Q0 nL0Q1 nL1Q0 VDD VSS PSRMND
XL1Q1 nL0Q2 nL0Q3 nL1Q1 VDD VSS PSRMND
XL1Q2 nL0Q4 nL0Q5 nL1Q2 VDD VSS PSRMND
XL1Q3 nL0Q6 nL0Q7 nL1Q3 VDD VSS PSRMND
XL1Q4 nL0Q8 nL0Q9 nL1Q4 VDD VSS PSRMND
XL1Q5 nL0Q10 nL0Q11 nL1Q5 VDD VSS PSRMND
XL1Q6 nL0Q12 nL0Q13 nL1Q6 VDD VSS PSRMND
XL1Q7 nL0Q14 nL0Q15 nL1Q7 VDD VSS PSRMND
XL1Q8 nL0Q16 nL0Q17 nL1Q8 VDD VSS PSRMND
XL1Q9 nL0Q18 nL0Q19 nL1Q9 VDD VSS PSRMND
XL1Q10 nL0Q20 nL0Q21 nL1Q10 VDD VSS PSRMND
XL1Q11 nL0Q22 nL0Q23 nL1Q11 VDD VSS PSRMND
XL1Q12 nL0Q24 nL0Q25 nL1Q12 VDD VSS PSRMND
XL1Q13 nL0Q26 nL0Q27 nL1Q13 VDD VSS PSRMND
XL1Q14 nL0Q28 nL0Q29 nL1Q14 VDD VSS PSRMND
XL1Q15 nL0Q30 nL0Q31 nL1Q15 VDD VSS PSRMND
XL2Q0 nL1Q0 nL1Q1 nL2Q0 VDD VSS PSRMNR
XL2Q1 nL1Q2 nL1Q3 nL2Q1 VDD VSS PSRMNR
XL2Q2 nL1Q4 nL1Q5 nL2Q2 VDD VSS PSRMNR
XL2Q3 nL1Q6 nL1Q7 nL2Q3 VDD VSS PSRMNR
XL2Q4 nL1Q8 nL1Q9 nL2Q4 VDD VSS PSRMNR
XL2Q5 nL1Q10 nL1Q11 nL2Q5 VDD VSS PSRMNR
XL2Q6 nL1Q12 nL1Q13 nL2Q6 VDD VSS PSRMNR
XL2Q7 nL1Q14 nL1Q15 nL2Q7 VDD VSS PSRMNR
XL3Q0 nL2Q0 nL2Q1 nL3Q0 VDD VSS PSRMND
XL3Q1 nL2Q2 nL2Q3 nL3Q1 VDD VSS PSRMND
XL3Q2 nL2Q4 nL2Q5 nL3Q2 VDD VSS PSRMND
XL3Q3 nL2Q6 nL2Q7 nL3Q3 VDD VSS PSRMND
XL4Q0 nL3Q0 nL3Q1 nL4Q0 VDD VSS PSRMNR
XL4Q1 nL3Q2 nL3Q3 nL4Q1 VDD VSS PSRMNR
XL5Q0 nL4Q0 nL4Q1 nQ VDD VSS PSRMND
.ENDS

.SUBCKT PS32X32 CK RE RA0 RA1 RA2 RA3 RA4 RD0 RD1 RD2 RD3 RD4 RD5 RD6 RD7 RD8 RD9 RD10 RD11 RD12 RD13 RD14 RD15 RD16 RD17 RD18 RD19 RD20 RD21 RD22 RD23 RD24 RD25 RD26 RD27 RD28 RD29 RD30 RD31 WE WA0 WA1 WA2 WA3 WA4 WD0 WD1 WD2 WD3 WD4 WD5 WD6 WD7 WD8 WD9 WD10 WD11 WD12 WD13 WD14 WD15 WD16 WD17 WD18 WD19 WD20 WD21 WD22 WD23 WD24 WD25 WD26 WD27 WD28 WD29 WD30 WD31 VDD VSS
XRWCKG RE WE CK nRCKP nRCKN nWCKP nWCKN VDD VSS PSRWCKG
XAD nWCKP nWCKN nRA0 nRA1 nRA2 nRA3 nRA4 WA0 WA1 WA2 WA3 WA4 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 VDD VSS PSAD32
XWDREG0 WD0 nWCKP nWCKN nWD0 iw0 VDD VSS PSREG
XWDREG1 WD1 nWCKP nWCKN nWD1 iw1 VDD VSS PSREG
XWDREG2 WD2 nWCKP nWCKN nWD2 iw2 VDD VSS PSREG
XWDREG3 WD3 nWCKP nWCKN nWD3 iw3 VDD VSS PSREG
XWDREG4 WD4 nWCKP nWCKN nWD4 iw4 VDD VSS PSREG
XWDREG5 WD5 nWCKP nWCKN nWD5 iw5 VDD VSS PSREG
XWDREG6 WD6 nWCKP nWCKN nWD6 iw6 VDD VSS PSREG
XWDREG7 WD7 nWCKP nWCKN nWD7 iw7 VDD VSS PSREG
XWDREG8 WD8 nWCKP nWCKN nWD8 iw8 VDD VSS PSREG
XWDREG9 WD9 nWCKP nWCKN nWD9 iw9 VDD VSS PSREG
XWDREG10 WD10 nWCKP nWCKN nWD10 iw10 VDD VSS PSREG
XWDREG11 WD11 nWCKP nWCKN nWD11 iw11 VDD VSS PSREG
XWDREG12 WD12 nWCKP nWCKN nWD12 iw12 VDD VSS PSREG
XWDREG13 WD13 nWCKP nWCKN nWD13 iw13 VDD VSS PSREG
XWDREG14 WD14 nWCKP nWCKN nWD14 iw14 VDD VSS PSREG
XWDREG15 WD15 nWCKP nWCKN nWD15 iw15 VDD VSS PSREG
XWDREG16 WD16 nWCKP nWCKN nWD16 iw16 VDD VSS PSREG
XWDREG17 WD17 nWCKP nWCKN nWD17 iw17 VDD VSS PSREG
XWDREG18 WD18 nWCKP nWCKN nWD18 iw18 VDD VSS PSREG
XWDREG19 WD19 nWCKP nWCKN nWD19 iw19 VDD VSS PSREG
XWDREG20 WD20 nWCKP nWCKN nWD20 iw20 VDD VSS PSREG
XWDREG21 WD21 nWCKP nWCKN nWD21 iw21 VDD VSS PSREG
XWDREG22 WD22 nWCKP nWCKN nWD22 iw22 VDD VSS PSREG
XWDREG23 WD23 nWCKP nWCKN nWD23 iw23 VDD VSS PSREG
XWDREG24 WD24 nWCKP nWCKN nWD24 iw24 VDD VSS PSREG
XWDREG25 WD25 nWCKP nWCKN nWD25 iw25 VDD VSS PSREG
XWDREG26 WD26 nWCKP nWCKN nWD26 iw26 VDD VSS PSREG
XWDREG27 WD27 nWCKP nWCKN nWD27 iw27 VDD VSS PSREG
XWDREG28 WD28 nWCKP nWCKN nWD28 iw28 VDD VSS PSREG
XWDREG29 WD29 nWCKP nWCKN nWD29 iw29 VDD VSS PSREG
XWDREG30 WD30 nWCKP nWCKN nWD30 iw30 VDD VSS PSREG
XWDREG31 WD31 nWCKP nWCKN nWD31 iw31 VDD VSS PSREG
XRAREG0 RA0 nRCKP nRCKN nRA0 ir0 VDD VSS PSREG
XRAREG1 RA1 nRCKP nRCKN nRA1 ir1 VDD VSS PSREG
XRAREG2 RA2 nRCKP nRCKN nRA2 ir2 VDD VSS PSREG
XRAREG3 RA3 nRCKP nRCKN nRA3 ir3 VDD VSS PSREG
XRAREG4 RA4 nRCKP nRCKN nRA4 ir4 VDD VSS PSREG
XBA0 nWD0 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD0 VDD VSS PSBA32
XBA1 nWD1 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD1 VDD VSS PSBA32
XBA2 nWD2 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD2 VDD VSS PSBA32
XBA3 nWD3 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD3 VDD VSS PSBA32
XBA4 nWD4 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD4 VDD VSS PSBA32
XBA5 nWD5 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD5 VDD VSS PSBA32
XBA6 nWD6 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD6 VDD VSS PSBA32
XBA7 nWD7 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD7 VDD VSS PSBA32
XBA8 nWD8 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD8 VDD VSS PSBA32
XBA9 nWD9 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD9 VDD VSS PSBA32
XBA10 nWD10 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD10 VDD VSS PSBA32
XBA11 nWD11 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD11 VDD VSS PSBA32
XBA12 nWD12 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD12 VDD VSS PSBA32
XBA13 nWD13 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD13 VDD VSS PSBA32
XBA14 nWD14 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD14 VDD VSS PSBA32
XBA15 nWD15 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD15 VDD VSS PSBA32
XBA16 nWD16 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD16 VDD VSS PSBA32
XBA17 nWD17 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD17 VDD VSS PSBA32
XBA18 nWD18 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD18 VDD VSS PSBA32
XBA19 nWD19 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD19 VDD VSS PSBA32
XBA20 nWD20 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD20 VDD VSS PSBA32
XBA21 nWD21 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD21 VDD VSS PSBA32
XBA22 nWD22 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD22 VDD VSS PSBA32
XBA23 nWD23 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD23 VDD VSS PSBA32
XBA24 nWD24 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD24 VDD VSS PSBA32
XBA25 nWD25 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD25 VDD VSS PSBA32
XBA26 nWD26 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD26 VDD VSS PSBA32
XBA27 nWD27 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD27 VDD VSS PSBA32
XBA28 nWD28 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD28 VDD VSS PSBA32
XBA29 nWD29 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD29 VDD VSS PSBA32
XBA30 nWD30 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD30 VDD VSS PSBA32
XBA31 nWD31 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 nS4 nGP4 nGN4 nS5 nGP5 nGN5 nS6 nGP6 nGN6 nS7 nGP7 nGN7 nS8 nGP8 nGN8 nS9 nGP9 nGN9 nS10 nGP10 nGN10 nS11 nGP11 nGN11 nS12 nGP12 nGN12 nS13 nGP13 nGN13 nS14 nGP14 nGN14 nS15 nGP15 nGN15 nS16 nGP16 nGN16 nS17 nGP17 nGN17 nS18 nGP18 nGN18 nS19 nGP19 nGN19 nS20 nGP20 nGN20 nS21 nGP21 nGN21 nS22 nGP22 nGN22 nS23 nGP23 nGN23 nS24 nGP24 nGN24 nS25 nGP25 nGN25 nS26 nGP26 nGN26 nS27 nGP27 nGN27 nS28 nGP28 nGN28 nS29 nGP29 nGN29 nS30 nGP30 nGN30 nS31 nGP31 nGN31 RD31 VDD VSS PSBA32
.ENDS
