.SUBCKT PSADOH4R A0 A1 Z VDD VSS
*.PININFO A0:I A1:I Z:O VDD:B VSS:B
X0 A0 A1 Z VDD VSS PSADOH_NR2
.ENDS

.SUBCKT PSADOH4 A0 A1 Z0 Z1 Z2 Z3 VDD VSS
XI0 A0 N0 VDD VSS PSADINV
XI1 A1 N1 VDD VSS PSADINV
X0 A0 A1 Z0 VDD VSS PSADOH4R
X1 N0 A1 Z1 VDD VSS PSADOH4R
X2 A0 N1 Z2 VDD VSS PSADOH4R
X3 N0 N1 Z3 VDD VSS PSADOH4R
.ENDS
