.SUBCKT PSBA4 D S0 GP0 GN0 S1 GP1 GN1 S2 GP2 GN2 S3 GP3 GN3 Q VDD VSS
X0 D GP0 GN0 S0 nL0Q0 VDD VSS PSBA1
X1 D GP1 GN1 S1 nL0Q1 VDD VSS PSBA1
X2 D GP2 GN2 S2 nL0Q2 VDD VSS PSBA1
X3 D GP3 GN3 S3 nL0Q3 VDD VSS PSBA1
XINV nQ Q VDD VSS PSRMINV
XL1Q0 nL0Q0 nL0Q1 nL1Q0 VDD VSS PSRMND
XL1Q1 nL0Q2 nL0Q3 nL1Q1 VDD VSS PSRMND
XL2Q0 nL1Q0 nL1Q1 nQ VDD VSS PSRMNR
.ENDS
