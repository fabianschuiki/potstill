.SUBCKT PSRMINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=450n L=60n M=1
.ENDS

.SUBCKT PSRMBUF A Z VDD VSS
MPM0 n1 A VDD VDD P_12_LLRVT W=210n L=60n M=1
MNM0 n1 A VSS VSS N_12_LLRVT W=150n L=60n M=1
MPM1 Z n1 VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM1 Z n1 VSS VSS N_12_LLRVT W=450n L=60n M=1
.ENDS

.SUBCKT PSRMND A B Z VDD VSS
*.PININFO A:I B:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=270n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=270n L=60n M=1
MNM0 Z B n1 VSS N_12_LLRVT W=180n L=60n M=1
MNM1 n1 A VSS VSS N_12_LLRVT W=180n L=60n M=1
.ENDS

.SUBCKT PSRMNR A B Z VDD VSS
*.PININFO A:I B:I Z:O
MPM0 n1 A VDD VDD P_12_LLRVT W=270n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=270n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=180n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=180n L=60n M=1
.ENDS

.SUBCKT PSADOH_ND2 A B Z VDD VSS
*.PININFO A:I B:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z B n1 VSS N_12_LLRVT W=480n L=60n M=1
MNM1 n1 A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_ND3 A B C Z VDD VSS
*.PININFO A:I B:I C:I Z:O VDD:B VSS:B
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM2 Z C VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z C n1 VSS N_12_LLRVT W=480n L=60n M=1
MNM1 n1 B n2 VSS N_12_LLRVT W=480n L=60n M=1
MNM2 n2 A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_NR2 A B Z VDD VSS
*.PININFO A:I B:I Z:O
MPM0 n1 A VDD VDD P_12_LLRVT W=660n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSADOH_NR3 A B C Z VDD VSS
*.PININFO A:I B:I C:I Z:O VDD:B VSS:B
MPM0 Z  C n1  VDD P_12_LLRVT W=660n L=60n M=1
MPM1 n1 B n2  VDD P_12_LLRVT W=660n L=60n M=1
MPM2 n2 A VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z  A VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM1 Z  B VSS VSS N_12_LLRVT W=480n L=60n M=1
MNM2 Z  C VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSREG_LA1 D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSREG_LA2 D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=300n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=450n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSREG D CKP CKN QP QN VDD VSS
XI0 D CKN CKP n1 i1 VDD VSS PSREG_LA1
XI1 n1 CKP CKN QP QN VDD VSS PSREG_LA2
.ENDS

.SUBCKT PSADCKG_LA D GP GN QP QN VDD VSS
MNM3 QP GN n1 VSS N_12_LLRVT W=150n L=60n M=1
MNM2 QP QN VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 QN n1 VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM0 D GP n1 VSS N_12_LLRVT W=150n L=60n M=1
MPM3 QP GP n1 VDD P_12_LLRVT W=150n L=60n M=1
MPM2 QP QN VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM1 QN n1 VDD VDD P_12_LLRVT W=150n L=60n M=1
MPM0 D GN n1 VDD P_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSADCKG_NR2 A B Z VDD VSS
MPM0 n1 A VDD VDD P_12_LLRVT W=630n L=60n M=1
MPM1 Z B n1 VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=150n L=60n M=1
MNM1 Z B VSS VSS N_12_LLRVT W=150n L=60n M=1
.ENDS

.SUBCKT PSADCKG E CKP CKN GCKP GCKN VDD VSS
X1 E CKN CKP i1 n1 VDD VSS PSADCKG_LA
X2 n1 CKN n2 VDD VSS PSADCKG_NR2
MPM0 GCKN n2 VDD VDD P_12_LLRVT W=600n L=60n M=1
MNM0 GCKN n2 VSS VSS N_12_LLRVT W=300n L=60n M=1
MPM1 GCKP GCKN VDD VDD P_12_LLRVT W=600n L=60n M=1
MNM1 GCKP GCKN VSS VSS N_12_LLRVT W=300n L=60n M=1
.ENDS

.SUBCKT PSADINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=660n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=480n L=60n M=1
.ENDS

.SUBCKT PSBA1 D GP GN S Q VDD VSS
*.PININFO D:I GP:I GN:I S:I Q:O VDD:B VSS:B
MNM0 net41 D VSS VSS N_12_LLRVT W=200e-9 L=60n M=1
MNM1 nFB GP net41 VSS N_12_LLRVT W=200e-9 L=60n M=1
MNM2 net40 nZ VSS VSS N_12_LLRVT W=150e-9 L=60n M=1
MNM3 nFB GN net40 VSS N_12_LLRVT W=150e-9 L=60n M=1
MNM4 nZ nFB VSS VSS N_12_LLRVT W=180e-9 L=60n M=1
MNM5 net42 S VSS VSS N_12_LLRVT W=180e-9 L=60n M=1
MNM6 Q nZ net42 VSS N_12_LLRVT W=180e-9 L=60n M=1
MPM0 nFB GN net38 VDD P_12_LLRVT W=300e-9 L=60n M=1
MPM1 net38 D VDD VDD P_12_LLRVT W=300e-9 L=60n M=1
MPM2 nFB GP net39 VDD P_12_LLRVT W=150e-9 L=60n M=1
MPM3 net39 nZ VDD VDD P_12_LLRVT W=150e-9 L=60n M=1
MPM4 nZ nFB VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
MPM5 Q nZ VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
MPM6 Q S VDD VDD P_12_LLRVT W=270e-9 L=60n M=1
.ENDS

.SUBCKT PSRWCKG_CKINV A Z VDD VSS
MPM0 Z A VDD VDD P_12_LLRVT W=630n L=60n M=1
MNM0 Z A VSS VSS N_12_LLRVT W=260n L=60n M=1
.ENDS

.SUBCKT PSRWCKG RE WE CK RCKP RCKN WCKP WCKN VDD VSS
X0 RE nCKP nCKN RCKP RCKN VDD VSS PSADCKG
X1 WE nCKP nCKN WCKP WCKN VDD VSS PSADCKG
X2 CK nCKN VDD VSS PSRWCKG_CKINV
X3 nCKN nCKP VDD VSS PSRWCKG_CKINV
.ENDS


.SUBCKT PSADOH4R A0 A1 Z VDD VSS
*.PININFO A0:I A1:I Z:O VDD:B VSS:B
X0 A0 A1 Z VDD VSS PSADOH_NR2
.ENDS

.SUBCKT PSADOH4 A0 A1 Z0 Z1 Z2 Z3 VDD VSS
XI0 A0 N0 VDD VSS PSADINV
XI1 A1 N1 VDD VSS PSADINV
X0 A0 A1 Z0 VDD VSS PSADOH4R
X1 N0 A1 Z1 VDD VSS PSADOH4R
X2 A0 N1 Z2 VDD VSS PSADOH4R
X3 N0 N1 Z3 VDD VSS PSADOH4R
.ENDS

.SUBCKT PSAD4 CKP CKN RA0 RA1 WA0 WA1 S0 GP0 GN0 S1 GP1 GN1 S2 GP2 GN2 S3 GP3 GN3 VDD VSS
XCKG0 nWE0 CKP CKN GP0 GN0 VDD VSS PSADCKG 
XCKG1 nWE1 CKP CKN GP1 GN1 VDD VSS PSADCKG 
XCKG2 nWE2 CKP CKN GP2 GN2 VDD VSS PSADCKG 
XCKG3 nWE3 CKP CKN GP3 GN3 VDD VSS PSADCKG 
XRAD RA0 RA1 S0 S1 S2 S3 VDD VSS PSADOH4
XWAD WA0 WA1 nWE0 nWE1 nWE2 nWE3 VDD VSS PSADOH4
.ENDS

.SUBCKT PSBA4 D S0 GP0 GN0 S1 GP1 GN1 S2 GP2 GN2 S3 GP3 GN3 Q VDD VSS
X0 D GP0 GN0 S0 nL0Q0 VDD VSS PSBA1
X1 D GP1 GN1 S1 nL0Q1 VDD VSS PSBA1
X2 D GP2 GN2 S2 nL0Q2 VDD VSS PSBA1
X3 D GP3 GN3 S3 nL0Q3 VDD VSS PSBA1
XINV nQ Q VDD VSS PSRMINV
XL1Q0 nL0Q0 nL0Q1 nL1Q0 VDD VSS PSRMND
XL1Q1 nL0Q2 nL0Q3 nL1Q1 VDD VSS PSRMND
XL2Q0 nL1Q0 nL1Q1 nQ VDD VSS PSRMNR
.ENDS

.SUBCKT PS4X128 CK RE RA0 RA1 RD0 RD1 RD2 RD3 RD4 RD5 RD6 RD7 RD8 RD9 RD10 RD11 RD12 RD13 RD14 RD15 RD16 RD17 RD18 RD19 RD20 RD21 RD22 RD23 RD24 RD25 RD26 RD27 RD28 RD29 RD30 RD31 RD32 RD33 RD34 RD35 RD36 RD37 RD38 RD39 RD40 RD41 RD42 RD43 RD44 RD45 RD46 RD47 RD48 RD49 RD50 RD51 RD52 RD53 RD54 RD55 RD56 RD57 RD58 RD59 RD60 RD61 RD62 RD63 RD64 RD65 RD66 RD67 RD68 RD69 RD70 RD71 RD72 RD73 RD74 RD75 RD76 RD77 RD78 RD79 RD80 RD81 RD82 RD83 RD84 RD85 RD86 RD87 RD88 RD89 RD90 RD91 RD92 RD93 RD94 RD95 RD96 RD97 RD98 RD99 RD100 RD101 RD102 RD103 RD104 RD105 RD106 RD107 RD108 RD109 RD110 RD111 RD112 RD113 RD114 RD115 RD116 RD117 RD118 RD119 RD120 RD121 RD122 RD123 RD124 RD125 RD126 RD127 WE WA0 WA1 WD0 WD1 WD2 WD3 WD4 WD5 WD6 WD7 WD8 WD9 WD10 WD11 WD12 WD13 WD14 WD15 WD16 WD17 WD18 WD19 WD20 WD21 WD22 WD23 WD24 WD25 WD26 WD27 WD28 WD29 WD30 WD31 WD32 WD33 WD34 WD35 WD36 WD37 WD38 WD39 WD40 WD41 WD42 WD43 WD44 WD45 WD46 WD47 WD48 WD49 WD50 WD51 WD52 WD53 WD54 WD55 WD56 WD57 WD58 WD59 WD60 WD61 WD62 WD63 WD64 WD65 WD66 WD67 WD68 WD69 WD70 WD71 WD72 WD73 WD74 WD75 WD76 WD77 WD78 WD79 WD80 WD81 WD82 WD83 WD84 WD85 WD86 WD87 WD88 WD89 WD90 WD91 WD92 WD93 WD94 WD95 WD96 WD97 WD98 WD99 WD100 WD101 WD102 WD103 WD104 WD105 WD106 WD107 WD108 WD109 WD110 WD111 WD112 WD113 WD114 WD115 WD116 WD117 WD118 WD119 WD120 WD121 WD122 WD123 WD124 WD125 WD126 WD127 VDD VSS
XRWCKG RE WE CK nRCKP nRCKN nWCKP nWCKN VDD VSS PSRWCKG
XAD nWCKP nWCKN nRA0 nRA1 WA0 WA1 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 VDD VSS PSAD4
XWDREG0 WD0 nWCKP nWCKN nWD0 iw0 VDD VSS PSREG
XWDREG1 WD1 nWCKP nWCKN nWD1 iw1 VDD VSS PSREG
XWDREG2 WD2 nWCKP nWCKN nWD2 iw2 VDD VSS PSREG
XWDREG3 WD3 nWCKP nWCKN nWD3 iw3 VDD VSS PSREG
XWDREG4 WD4 nWCKP nWCKN nWD4 iw4 VDD VSS PSREG
XWDREG5 WD5 nWCKP nWCKN nWD5 iw5 VDD VSS PSREG
XWDREG6 WD6 nWCKP nWCKN nWD6 iw6 VDD VSS PSREG
XWDREG7 WD7 nWCKP nWCKN nWD7 iw7 VDD VSS PSREG
XWDREG8 WD8 nWCKP nWCKN nWD8 iw8 VDD VSS PSREG
XWDREG9 WD9 nWCKP nWCKN nWD9 iw9 VDD VSS PSREG
XWDREG10 WD10 nWCKP nWCKN nWD10 iw10 VDD VSS PSREG
XWDREG11 WD11 nWCKP nWCKN nWD11 iw11 VDD VSS PSREG
XWDREG12 WD12 nWCKP nWCKN nWD12 iw12 VDD VSS PSREG
XWDREG13 WD13 nWCKP nWCKN nWD13 iw13 VDD VSS PSREG
XWDREG14 WD14 nWCKP nWCKN nWD14 iw14 VDD VSS PSREG
XWDREG15 WD15 nWCKP nWCKN nWD15 iw15 VDD VSS PSREG
XWDREG16 WD16 nWCKP nWCKN nWD16 iw16 VDD VSS PSREG
XWDREG17 WD17 nWCKP nWCKN nWD17 iw17 VDD VSS PSREG
XWDREG18 WD18 nWCKP nWCKN nWD18 iw18 VDD VSS PSREG
XWDREG19 WD19 nWCKP nWCKN nWD19 iw19 VDD VSS PSREG
XWDREG20 WD20 nWCKP nWCKN nWD20 iw20 VDD VSS PSREG
XWDREG21 WD21 nWCKP nWCKN nWD21 iw21 VDD VSS PSREG
XWDREG22 WD22 nWCKP nWCKN nWD22 iw22 VDD VSS PSREG
XWDREG23 WD23 nWCKP nWCKN nWD23 iw23 VDD VSS PSREG
XWDREG24 WD24 nWCKP nWCKN nWD24 iw24 VDD VSS PSREG
XWDREG25 WD25 nWCKP nWCKN nWD25 iw25 VDD VSS PSREG
XWDREG26 WD26 nWCKP nWCKN nWD26 iw26 VDD VSS PSREG
XWDREG27 WD27 nWCKP nWCKN nWD27 iw27 VDD VSS PSREG
XWDREG28 WD28 nWCKP nWCKN nWD28 iw28 VDD VSS PSREG
XWDREG29 WD29 nWCKP nWCKN nWD29 iw29 VDD VSS PSREG
XWDREG30 WD30 nWCKP nWCKN nWD30 iw30 VDD VSS PSREG
XWDREG31 WD31 nWCKP nWCKN nWD31 iw31 VDD VSS PSREG
XWDREG32 WD32 nWCKP nWCKN nWD32 iw32 VDD VSS PSREG
XWDREG33 WD33 nWCKP nWCKN nWD33 iw33 VDD VSS PSREG
XWDREG34 WD34 nWCKP nWCKN nWD34 iw34 VDD VSS PSREG
XWDREG35 WD35 nWCKP nWCKN nWD35 iw35 VDD VSS PSREG
XWDREG36 WD36 nWCKP nWCKN nWD36 iw36 VDD VSS PSREG
XWDREG37 WD37 nWCKP nWCKN nWD37 iw37 VDD VSS PSREG
XWDREG38 WD38 nWCKP nWCKN nWD38 iw38 VDD VSS PSREG
XWDREG39 WD39 nWCKP nWCKN nWD39 iw39 VDD VSS PSREG
XWDREG40 WD40 nWCKP nWCKN nWD40 iw40 VDD VSS PSREG
XWDREG41 WD41 nWCKP nWCKN nWD41 iw41 VDD VSS PSREG
XWDREG42 WD42 nWCKP nWCKN nWD42 iw42 VDD VSS PSREG
XWDREG43 WD43 nWCKP nWCKN nWD43 iw43 VDD VSS PSREG
XWDREG44 WD44 nWCKP nWCKN nWD44 iw44 VDD VSS PSREG
XWDREG45 WD45 nWCKP nWCKN nWD45 iw45 VDD VSS PSREG
XWDREG46 WD46 nWCKP nWCKN nWD46 iw46 VDD VSS PSREG
XWDREG47 WD47 nWCKP nWCKN nWD47 iw47 VDD VSS PSREG
XWDREG48 WD48 nWCKP nWCKN nWD48 iw48 VDD VSS PSREG
XWDREG49 WD49 nWCKP nWCKN nWD49 iw49 VDD VSS PSREG
XWDREG50 WD50 nWCKP nWCKN nWD50 iw50 VDD VSS PSREG
XWDREG51 WD51 nWCKP nWCKN nWD51 iw51 VDD VSS PSREG
XWDREG52 WD52 nWCKP nWCKN nWD52 iw52 VDD VSS PSREG
XWDREG53 WD53 nWCKP nWCKN nWD53 iw53 VDD VSS PSREG
XWDREG54 WD54 nWCKP nWCKN nWD54 iw54 VDD VSS PSREG
XWDREG55 WD55 nWCKP nWCKN nWD55 iw55 VDD VSS PSREG
XWDREG56 WD56 nWCKP nWCKN nWD56 iw56 VDD VSS PSREG
XWDREG57 WD57 nWCKP nWCKN nWD57 iw57 VDD VSS PSREG
XWDREG58 WD58 nWCKP nWCKN nWD58 iw58 VDD VSS PSREG
XWDREG59 WD59 nWCKP nWCKN nWD59 iw59 VDD VSS PSREG
XWDREG60 WD60 nWCKP nWCKN nWD60 iw60 VDD VSS PSREG
XWDREG61 WD61 nWCKP nWCKN nWD61 iw61 VDD VSS PSREG
XWDREG62 WD62 nWCKP nWCKN nWD62 iw62 VDD VSS PSREG
XWDREG63 WD63 nWCKP nWCKN nWD63 iw63 VDD VSS PSREG
XWDREG64 WD64 nWCKP nWCKN nWD64 iw64 VDD VSS PSREG
XWDREG65 WD65 nWCKP nWCKN nWD65 iw65 VDD VSS PSREG
XWDREG66 WD66 nWCKP nWCKN nWD66 iw66 VDD VSS PSREG
XWDREG67 WD67 nWCKP nWCKN nWD67 iw67 VDD VSS PSREG
XWDREG68 WD68 nWCKP nWCKN nWD68 iw68 VDD VSS PSREG
XWDREG69 WD69 nWCKP nWCKN nWD69 iw69 VDD VSS PSREG
XWDREG70 WD70 nWCKP nWCKN nWD70 iw70 VDD VSS PSREG
XWDREG71 WD71 nWCKP nWCKN nWD71 iw71 VDD VSS PSREG
XWDREG72 WD72 nWCKP nWCKN nWD72 iw72 VDD VSS PSREG
XWDREG73 WD73 nWCKP nWCKN nWD73 iw73 VDD VSS PSREG
XWDREG74 WD74 nWCKP nWCKN nWD74 iw74 VDD VSS PSREG
XWDREG75 WD75 nWCKP nWCKN nWD75 iw75 VDD VSS PSREG
XWDREG76 WD76 nWCKP nWCKN nWD76 iw76 VDD VSS PSREG
XWDREG77 WD77 nWCKP nWCKN nWD77 iw77 VDD VSS PSREG
XWDREG78 WD78 nWCKP nWCKN nWD78 iw78 VDD VSS PSREG
XWDREG79 WD79 nWCKP nWCKN nWD79 iw79 VDD VSS PSREG
XWDREG80 WD80 nWCKP nWCKN nWD80 iw80 VDD VSS PSREG
XWDREG81 WD81 nWCKP nWCKN nWD81 iw81 VDD VSS PSREG
XWDREG82 WD82 nWCKP nWCKN nWD82 iw82 VDD VSS PSREG
XWDREG83 WD83 nWCKP nWCKN nWD83 iw83 VDD VSS PSREG
XWDREG84 WD84 nWCKP nWCKN nWD84 iw84 VDD VSS PSREG
XWDREG85 WD85 nWCKP nWCKN nWD85 iw85 VDD VSS PSREG
XWDREG86 WD86 nWCKP nWCKN nWD86 iw86 VDD VSS PSREG
XWDREG87 WD87 nWCKP nWCKN nWD87 iw87 VDD VSS PSREG
XWDREG88 WD88 nWCKP nWCKN nWD88 iw88 VDD VSS PSREG
XWDREG89 WD89 nWCKP nWCKN nWD89 iw89 VDD VSS PSREG
XWDREG90 WD90 nWCKP nWCKN nWD90 iw90 VDD VSS PSREG
XWDREG91 WD91 nWCKP nWCKN nWD91 iw91 VDD VSS PSREG
XWDREG92 WD92 nWCKP nWCKN nWD92 iw92 VDD VSS PSREG
XWDREG93 WD93 nWCKP nWCKN nWD93 iw93 VDD VSS PSREG
XWDREG94 WD94 nWCKP nWCKN nWD94 iw94 VDD VSS PSREG
XWDREG95 WD95 nWCKP nWCKN nWD95 iw95 VDD VSS PSREG
XWDREG96 WD96 nWCKP nWCKN nWD96 iw96 VDD VSS PSREG
XWDREG97 WD97 nWCKP nWCKN nWD97 iw97 VDD VSS PSREG
XWDREG98 WD98 nWCKP nWCKN nWD98 iw98 VDD VSS PSREG
XWDREG99 WD99 nWCKP nWCKN nWD99 iw99 VDD VSS PSREG
XWDREG100 WD100 nWCKP nWCKN nWD100 iw100 VDD VSS PSREG
XWDREG101 WD101 nWCKP nWCKN nWD101 iw101 VDD VSS PSREG
XWDREG102 WD102 nWCKP nWCKN nWD102 iw102 VDD VSS PSREG
XWDREG103 WD103 nWCKP nWCKN nWD103 iw103 VDD VSS PSREG
XWDREG104 WD104 nWCKP nWCKN nWD104 iw104 VDD VSS PSREG
XWDREG105 WD105 nWCKP nWCKN nWD105 iw105 VDD VSS PSREG
XWDREG106 WD106 nWCKP nWCKN nWD106 iw106 VDD VSS PSREG
XWDREG107 WD107 nWCKP nWCKN nWD107 iw107 VDD VSS PSREG
XWDREG108 WD108 nWCKP nWCKN nWD108 iw108 VDD VSS PSREG
XWDREG109 WD109 nWCKP nWCKN nWD109 iw109 VDD VSS PSREG
XWDREG110 WD110 nWCKP nWCKN nWD110 iw110 VDD VSS PSREG
XWDREG111 WD111 nWCKP nWCKN nWD111 iw111 VDD VSS PSREG
XWDREG112 WD112 nWCKP nWCKN nWD112 iw112 VDD VSS PSREG
XWDREG113 WD113 nWCKP nWCKN nWD113 iw113 VDD VSS PSREG
XWDREG114 WD114 nWCKP nWCKN nWD114 iw114 VDD VSS PSREG
XWDREG115 WD115 nWCKP nWCKN nWD115 iw115 VDD VSS PSREG
XWDREG116 WD116 nWCKP nWCKN nWD116 iw116 VDD VSS PSREG
XWDREG117 WD117 nWCKP nWCKN nWD117 iw117 VDD VSS PSREG
XWDREG118 WD118 nWCKP nWCKN nWD118 iw118 VDD VSS PSREG
XWDREG119 WD119 nWCKP nWCKN nWD119 iw119 VDD VSS PSREG
XWDREG120 WD120 nWCKP nWCKN nWD120 iw120 VDD VSS PSREG
XWDREG121 WD121 nWCKP nWCKN nWD121 iw121 VDD VSS PSREG
XWDREG122 WD122 nWCKP nWCKN nWD122 iw122 VDD VSS PSREG
XWDREG123 WD123 nWCKP nWCKN nWD123 iw123 VDD VSS PSREG
XWDREG124 WD124 nWCKP nWCKN nWD124 iw124 VDD VSS PSREG
XWDREG125 WD125 nWCKP nWCKN nWD125 iw125 VDD VSS PSREG
XWDREG126 WD126 nWCKP nWCKN nWD126 iw126 VDD VSS PSREG
XWDREG127 WD127 nWCKP nWCKN nWD127 iw127 VDD VSS PSREG
XRAREG0 RA0 nRCKP nRCKN nRA0 ir0 VDD VSS PSREG
XRAREG1 RA1 nRCKP nRCKN nRA1 ir1 VDD VSS PSREG
XBA0 nWD0 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD0 VDD VSS PSBA4
XBA1 nWD1 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD1 VDD VSS PSBA4
XBA2 nWD2 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD2 VDD VSS PSBA4
XBA3 nWD3 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD3 VDD VSS PSBA4
XBA4 nWD4 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD4 VDD VSS PSBA4
XBA5 nWD5 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD5 VDD VSS PSBA4
XBA6 nWD6 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD6 VDD VSS PSBA4
XBA7 nWD7 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD7 VDD VSS PSBA4
XBA8 nWD8 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD8 VDD VSS PSBA4
XBA9 nWD9 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD9 VDD VSS PSBA4
XBA10 nWD10 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD10 VDD VSS PSBA4
XBA11 nWD11 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD11 VDD VSS PSBA4
XBA12 nWD12 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD12 VDD VSS PSBA4
XBA13 nWD13 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD13 VDD VSS PSBA4
XBA14 nWD14 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD14 VDD VSS PSBA4
XBA15 nWD15 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD15 VDD VSS PSBA4
XBA16 nWD16 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD16 VDD VSS PSBA4
XBA17 nWD17 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD17 VDD VSS PSBA4
XBA18 nWD18 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD18 VDD VSS PSBA4
XBA19 nWD19 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD19 VDD VSS PSBA4
XBA20 nWD20 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD20 VDD VSS PSBA4
XBA21 nWD21 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD21 VDD VSS PSBA4
XBA22 nWD22 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD22 VDD VSS PSBA4
XBA23 nWD23 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD23 VDD VSS PSBA4
XBA24 nWD24 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD24 VDD VSS PSBA4
XBA25 nWD25 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD25 VDD VSS PSBA4
XBA26 nWD26 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD26 VDD VSS PSBA4
XBA27 nWD27 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD27 VDD VSS PSBA4
XBA28 nWD28 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD28 VDD VSS PSBA4
XBA29 nWD29 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD29 VDD VSS PSBA4
XBA30 nWD30 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD30 VDD VSS PSBA4
XBA31 nWD31 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD31 VDD VSS PSBA4
XBA32 nWD32 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD32 VDD VSS PSBA4
XBA33 nWD33 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD33 VDD VSS PSBA4
XBA34 nWD34 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD34 VDD VSS PSBA4
XBA35 nWD35 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD35 VDD VSS PSBA4
XBA36 nWD36 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD36 VDD VSS PSBA4
XBA37 nWD37 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD37 VDD VSS PSBA4
XBA38 nWD38 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD38 VDD VSS PSBA4
XBA39 nWD39 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD39 VDD VSS PSBA4
XBA40 nWD40 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD40 VDD VSS PSBA4
XBA41 nWD41 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD41 VDD VSS PSBA4
XBA42 nWD42 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD42 VDD VSS PSBA4
XBA43 nWD43 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD43 VDD VSS PSBA4
XBA44 nWD44 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD44 VDD VSS PSBA4
XBA45 nWD45 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD45 VDD VSS PSBA4
XBA46 nWD46 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD46 VDD VSS PSBA4
XBA47 nWD47 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD47 VDD VSS PSBA4
XBA48 nWD48 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD48 VDD VSS PSBA4
XBA49 nWD49 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD49 VDD VSS PSBA4
XBA50 nWD50 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD50 VDD VSS PSBA4
XBA51 nWD51 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD51 VDD VSS PSBA4
XBA52 nWD52 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD52 VDD VSS PSBA4
XBA53 nWD53 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD53 VDD VSS PSBA4
XBA54 nWD54 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD54 VDD VSS PSBA4
XBA55 nWD55 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD55 VDD VSS PSBA4
XBA56 nWD56 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD56 VDD VSS PSBA4
XBA57 nWD57 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD57 VDD VSS PSBA4
XBA58 nWD58 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD58 VDD VSS PSBA4
XBA59 nWD59 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD59 VDD VSS PSBA4
XBA60 nWD60 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD60 VDD VSS PSBA4
XBA61 nWD61 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD61 VDD VSS PSBA4
XBA62 nWD62 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD62 VDD VSS PSBA4
XBA63 nWD63 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD63 VDD VSS PSBA4
XBA64 nWD64 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD64 VDD VSS PSBA4
XBA65 nWD65 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD65 VDD VSS PSBA4
XBA66 nWD66 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD66 VDD VSS PSBA4
XBA67 nWD67 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD67 VDD VSS PSBA4
XBA68 nWD68 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD68 VDD VSS PSBA4
XBA69 nWD69 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD69 VDD VSS PSBA4
XBA70 nWD70 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD70 VDD VSS PSBA4
XBA71 nWD71 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD71 VDD VSS PSBA4
XBA72 nWD72 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD72 VDD VSS PSBA4
XBA73 nWD73 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD73 VDD VSS PSBA4
XBA74 nWD74 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD74 VDD VSS PSBA4
XBA75 nWD75 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD75 VDD VSS PSBA4
XBA76 nWD76 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD76 VDD VSS PSBA4
XBA77 nWD77 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD77 VDD VSS PSBA4
XBA78 nWD78 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD78 VDD VSS PSBA4
XBA79 nWD79 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD79 VDD VSS PSBA4
XBA80 nWD80 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD80 VDD VSS PSBA4
XBA81 nWD81 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD81 VDD VSS PSBA4
XBA82 nWD82 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD82 VDD VSS PSBA4
XBA83 nWD83 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD83 VDD VSS PSBA4
XBA84 nWD84 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD84 VDD VSS PSBA4
XBA85 nWD85 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD85 VDD VSS PSBA4
XBA86 nWD86 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD86 VDD VSS PSBA4
XBA87 nWD87 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD87 VDD VSS PSBA4
XBA88 nWD88 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD88 VDD VSS PSBA4
XBA89 nWD89 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD89 VDD VSS PSBA4
XBA90 nWD90 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD90 VDD VSS PSBA4
XBA91 nWD91 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD91 VDD VSS PSBA4
XBA92 nWD92 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD92 VDD VSS PSBA4
XBA93 nWD93 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD93 VDD VSS PSBA4
XBA94 nWD94 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD94 VDD VSS PSBA4
XBA95 nWD95 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD95 VDD VSS PSBA4
XBA96 nWD96 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD96 VDD VSS PSBA4
XBA97 nWD97 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD97 VDD VSS PSBA4
XBA98 nWD98 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD98 VDD VSS PSBA4
XBA99 nWD99 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD99 VDD VSS PSBA4
XBA100 nWD100 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD100 VDD VSS PSBA4
XBA101 nWD101 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD101 VDD VSS PSBA4
XBA102 nWD102 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD102 VDD VSS PSBA4
XBA103 nWD103 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD103 VDD VSS PSBA4
XBA104 nWD104 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD104 VDD VSS PSBA4
XBA105 nWD105 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD105 VDD VSS PSBA4
XBA106 nWD106 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD106 VDD VSS PSBA4
XBA107 nWD107 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD107 VDD VSS PSBA4
XBA108 nWD108 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD108 VDD VSS PSBA4
XBA109 nWD109 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD109 VDD VSS PSBA4
XBA110 nWD110 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD110 VDD VSS PSBA4
XBA111 nWD111 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD111 VDD VSS PSBA4
XBA112 nWD112 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD112 VDD VSS PSBA4
XBA113 nWD113 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD113 VDD VSS PSBA4
XBA114 nWD114 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD114 VDD VSS PSBA4
XBA115 nWD115 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD115 VDD VSS PSBA4
XBA116 nWD116 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD116 VDD VSS PSBA4
XBA117 nWD117 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD117 VDD VSS PSBA4
XBA118 nWD118 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD118 VDD VSS PSBA4
XBA119 nWD119 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD119 VDD VSS PSBA4
XBA120 nWD120 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD120 VDD VSS PSBA4
XBA121 nWD121 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD121 VDD VSS PSBA4
XBA122 nWD122 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD122 VDD VSS PSBA4
XBA123 nWD123 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD123 VDD VSS PSBA4
XBA124 nWD124 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD124 VDD VSS PSBA4
XBA125 nWD125 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD125 VDD VSS PSBA4
XBA126 nWD126 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD126 VDD VSS PSBA4
XBA127 nWD127 nS0 nGP0 nGN0 nS1 nGP1 nGN1 nS2 nGP2 nGN2 nS3 nGP3 nGN3 RD127 VDD VSS PSBA4
.ENDS
