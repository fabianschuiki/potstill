.SUBCKT PSADOH4R A0 A1 Z VDD VSS
*.PININFO A0:I A1:I Z:O VDD:B VSS:B
X0 A0 A1 Z VDD VSS PSADOH_NR2
.ENDS

.SUBCKT PSADOH4 A0 A1 Z0 Z1 Z2 Z3 VDD VSS
XI0 A0 N0 VDD VSS PSADINV
XI1 A1 N1 VDD VSS PSADINV
X0 A0 A1 Z0 VDD VSS PSADOH4R
X1 N0 A1 Z1 VDD VSS PSADOH4R
X2 A0 N1 Z2 VDD VSS PSADOH4R
X3 N0 N1 Z3 VDD VSS PSADOH4R
.ENDS

.SUBCKT PSAD4 CKP CKN RA0 RA1 WA0 WA1 S0 GP0 GN0 S1 GP1 GN1 S2 GP2 GN2 S3 GP3 GN3 VDD VSS
XCKG0 nWE0 CKP CKN GP0 GN0 VDD VSS PSADCKG 
XCKG1 nWE1 CKP CKN GP1 GN1 VDD VSS PSADCKG 
XCKG2 nWE2 CKP CKN GP2 GN2 VDD VSS PSADCKG 
XCKG3 nWE3 CKP CKN GP3 GN3 VDD VSS PSADCKG 
XRAD RA0 RA1 S0 S1 S2 S3 VDD VSS PSADOH4
XWAD WA0 WA1 nWE0 nWE1 nWE2 nWE3 VDD VSS PSADOH4
.ENDS
